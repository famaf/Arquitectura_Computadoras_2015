library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity imem is
    port (
            a : in std_logic_vector (5 DOWNTO 0);
            y : out std_logic_vector (31 DOWNTO 0)
         );
end imem;


architecture memory of imem is

    type memoria_rom is array (0 to 63) of std_logic_vector (31 downto 0);

    signal myrom : memoria_rom := (
    "11110000000000000000000000000000", -- 00000000 -- 0
    "11110000000000000000000000000001", -- 00000001 -- 1
    "00000000000000000000000000000010", -- 00000002 -- 2
    "00000000000000000000000000000011", -- 00000003 -- 3
    "00000000000000000000000000000100", -- 00000004 -- 4
    "00000000000000000000000000000101", -- 00000005 -- 5
    "00000000000000000000000000000110", -- 00000006 -- 6
    "00000000000000000000000000000111", -- 00000007 -- 7
    "00000000000000000000000000001000", -- 00000008 -- 8
    "00000000000000000000000000001001", -- 00000009 -- 9
    "00000000000000000000000000001010", -- 0000000A -- 10
    "00000000000000000000000000001011", -- 0000000B -- 11
    "00000000000000000000000000001100", -- 0000000C -- 12
    "00000000000000000000000000001101", -- 0000000D -- 13
    "00000000000000000000000000001110", -- 0000000E -- 14
    "00000000000000000000000000001111", -- 0000000F -- 15
    "00000000000000000000000000010000", -- 00000010 -- 16
    "00000000000000000000000000010001", -- 00000011 -- 17 
    "00000000000000000000000000010010", -- 00000012 -- 18
    "00000000000000000000000000010011", -- 00000013 -- 19
    "00000000000000000000000000010100", -- 00000014 -- 20
    "00000000000000000000000000010101", -- 00000015 -- 21
    "00000000000000000000000000010110", -- 00000016 -- 22
    "00000000000000000000000000010111", -- 00000017 -- 23
    "00000000000000000000000000011000", -- 00000018 -- 24
    "00000000000000000000000000011001", -- 00000019 -- 25
    "00000000000000000000000000011010", -- 0000001A -- 26
    "00000000000000000000000000011011", -- 0000001B -- 27
    "00000000000000000000000000011100", -- 0000001C -- 28
    "00000000000000000000000000011101", -- 0000001D -- 29
    "00000000000000000000000000011110", -- 0000001E -- 30
    "00000000000000000000000000011111", -- 0000001F -- 31
    "00000000000000000000000000100000", -- 00000020 -- 32
    "00000000000000000000000000100001", -- 00000021 -- 33
    "00000000000000000000000000100010", -- 00000022 -- 34
    "00000000000000000000000000100011", -- 00000023 -- 35
    "00000000000000000000000000100100", -- 00000024 -- 36
    "00000000000000000000000000100101", -- 00000025 -- 37
    "00000000000000000000000000100110", -- 00000026 -- 38
    "00000000000000000000000000100111", -- 00000027 -- 39
    "00000000000000000000000000101000", -- 00000028 -- 40
    "00000000000000000000000000101001", -- 00000029 -- 41
    "00000000000000000000000000101010", -- 0000002A -- 42
    "00000000000000000000000000101011", -- 0000002B -- 43
    "00000000000000000000000000101100", -- 0000002C -- 44
    "00000000000000000000000000101101", -- 0000002D -- 45
    "00000000000000000000000000101110", -- 0000002E -- 46
    "00000000000000000000000000101111", -- 0000002F -- 47
    "00000000000000000000000000110000", -- 00000030 -- 48
    "00000000000000000000000000110001", -- 00000031 -- 49
    "00000000000000000000000000110010", -- 00000032 -- 50
    "00000000000000000000000000110011", -- 00000033 -- 51
    "00000000000000000000000000110100", -- 00000034 -- 52
    "00000000000000000000000000110101", -- 00000035 -- 53
    "00000000000000000000000000110110", -- 00000036 -- 54
    "00000000000000000000000000110111", -- 00000037 -- 55
    "00000000000000000000000000111000", -- 00000038 -- 56
    "00000000000000000000000000111001", -- 00000039 -- 57
    "00000000000000000000000000111010", -- 0000003A -- 58
    "00000000000000000000000000111011", -- 0000003B -- 59
    "00000000000000000000000000111100", -- 0000003C -- 60
    "00000000000000000000000000111101", -- 0000003D -- 61
    "00000000000000000000000000111110", -- 0000003E -- 62
    "11110000000000000000000000111111" -- 0000003F -- 63
    );

begin

    process (a) begin
        y <= myrom(to_integer(unsigned(a)));
    end process;
end memory;

-- VER WARNING AL COMPILAR
